/*

Any particular permutation of 8 digits from 1 to 8
can be produced by swapping (first number, another number)
10 times, for example

1 2 3 4 5 6 7 8
5 2 3 4 1 6 7 8
4 2 3 5 1 6 7 8
1 2 3 5 4 6 7 8
3 2 1 5 4 6 7 8
6 2 1 5 4 3 7 8
1 2 6 5 4 3 7 8
7 2 6 5 4 3 1 8
2 7 6 5 4 3 1 8
1 7 6 5 4 3 2 8
8 7 6 5 4 3 2 1

as such, the shift_key is ideally 10 x 3 bits in length.

However, we make do with 8 x 3 bits for now. 

*/

module GenPermutateKey (
    // input shift key
    input   wire [23:0] shift_key,
    // permute_key1 is for first 8 samples
    // permute_key2 is for last 8 samples
    // permute_key2 is reverse of permute_key1
    output  wire [23:0] permute_key1,
    output  wire [23:0] permute_key2
);

    wire [23:0] tmp0, tmp1, tmp2, tmp3, tmp4, tmp5, tmp6, tmp7;
    wire [2:0]  k0, k1, k2, k3, k4, k5, k6, k7; // for readability + debugging

// number  1
assign k0 = shift_key[23:21];
assign tmp0 =   (k0 == 'b000) ? {3'd0, 3'd1, 3'd2, 3'd3, 3'd4, 3'd5, 3'd6, 3'd7} :
                (k0 == 'b001) ? {3'd1, 3'd0, 3'd2, 3'd3, 3'd4, 3'd5, 3'd6, 3'd7} :
                (k0 == 'b010) ? {3'd2, 3'd1, 3'd0, 3'd3, 3'd4, 3'd5, 3'd6, 3'd7} :
                (k0 == 'b011) ? {3'd3, 3'd1, 3'd2, 3'd0, 3'd4, 3'd5, 3'd6, 3'd7} :
                (k0 == 'b100) ? {3'd4, 3'd1, 3'd2, 3'd3, 3'd0, 3'd5, 3'd6, 3'd7} :
                (k0 == 'b101) ? {3'd5, 3'd1, 3'd2, 3'd3, 3'd4, 3'd0, 3'd6, 3'd7} :
                (k0 == 'b110) ? {3'd6, 3'd1, 3'd2, 3'd3, 3'd4, 3'd5, 3'd0, 3'd7} :
                (k0 == 'b111) ? {3'd7, 3'd1, 3'd2, 3'd3, 3'd4, 3'd5, 3'd6, 3'd0} :
                                3'bx ;

// number 2
assign k1 = shift_key[20:18];
assign tmp1 =   (k1 == 'b000) ? {tmp0[23:21], tmp0[20:18], tmp0[17:15], tmp0[14:12], tmp0[11:09], tmp0[08:06], tmp0[05:03], tmp0[02:00]} :
                (k1 == 'b001) ? {tmp0[20:18], tmp0[23:21], tmp0[17:15], tmp0[14:12], tmp0[11:09], tmp0[08:06], tmp0[05:03], tmp0[02:00]} :
                (k1 == 'b010) ? {tmp0[17:15], tmp0[20:18], tmp0[23:21], tmp0[14:12], tmp0[11:09], tmp0[08:06], tmp0[05:03], tmp0[02:00]} :
                (k1 == 'b011) ? {tmp0[14:12], tmp0[20:18], tmp0[17:15], tmp0[23:21], tmp0[11:09], tmp0[08:06], tmp0[05:03], tmp0[02:00]} :
                (k1 == 'b100) ? {tmp0[11:09], tmp0[20:18], tmp0[17:15], tmp0[14:12], tmp0[23:21], tmp0[08:06], tmp0[05:03], tmp0[02:00]} :
                (k1 == 'b101) ? {tmp0[08:06], tmp0[20:18], tmp0[17:15], tmp0[14:12], tmp0[11:09], tmp0[23:21], tmp0[05:03], tmp0[02:00]} :
                (k1 == 'b110) ? {tmp0[05:03], tmp0[20:18], tmp0[17:15], tmp0[14:12], tmp0[11:09], tmp0[08:06], tmp0[23:21], tmp0[02:00]} :
                (k1 == 'b111) ? {tmp0[02:00], tmp0[20:18], tmp0[17:15], tmp0[14:12], tmp0[11:09], tmp0[08:06], tmp0[05:03], tmp0[23:21]} :
                                3'bx ;

// number 3
assign k2 = shift_key[17:15];
assign tmp2 =   (k2 == 'b000) ? {tmp1[23:21], tmp1[20:18], tmp1[17:15], tmp1[14:12], tmp1[11:09], tmp1[08:06], tmp1[05:03], tmp1[02:00]} :
                (k2 == 'b001) ? {tmp1[20:18], tmp1[23:21], tmp1[17:15], tmp1[14:12], tmp1[11:09], tmp1[08:06], tmp1[05:03], tmp1[02:00]} :
                (k2 == 'b010) ? {tmp1[17:15], tmp1[20:18], tmp1[23:21], tmp1[14:12], tmp1[11:09], tmp1[08:06], tmp1[05:03], tmp1[02:00]} :
                (k2 == 'b011) ? {tmp1[14:12], tmp1[20:18], tmp1[17:15], tmp1[23:21], tmp1[11:09], tmp1[08:06], tmp1[05:03], tmp1[02:00]} :
                (k2 == 'b100) ? {tmp1[11:09], tmp1[20:18], tmp1[17:15], tmp1[14:12], tmp1[23:21], tmp1[08:06], tmp1[05:03], tmp1[02:00]} :
                (k2 == 'b101) ? {tmp1[08:06], tmp1[20:18], tmp1[17:15], tmp1[14:12], tmp1[11:09], tmp1[23:21], tmp1[05:03], tmp1[02:00]} :
                (k2 == 'b110) ? {tmp1[05:03], tmp1[20:18], tmp1[17:15], tmp1[14:12], tmp1[11:09], tmp1[08:06], tmp1[23:21], tmp1[02:00]} :
                (k2 == 'b111) ? {tmp1[02:00], tmp1[20:18], tmp1[17:15], tmp1[14:12], tmp1[11:09], tmp1[08:06], tmp1[05:03], tmp1[23:21]} :
                                3'bx ;

// number 4
assign k3 = shift_key[14:12];
assign tmp3 =   (k3 == 'b000) ? {tmp2[23:21], tmp2[20:18], tmp2[17:15], tmp2[14:12], tmp2[11:09], tmp2[08:06], tmp2[05:03], tmp2[02:00]} :
                (k3 == 'b001) ? {tmp2[20:18], tmp2[23:21], tmp2[17:15], tmp2[14:12], tmp2[11:09], tmp2[08:06], tmp2[05:03], tmp2[02:00]} :
                (k3 == 'b010) ? {tmp2[17:15], tmp2[20:18], tmp2[23:21], tmp2[14:12], tmp2[11:09], tmp2[08:06], tmp2[05:03], tmp2[02:00]} :
                (k3 == 'b011) ? {tmp2[14:12], tmp2[20:18], tmp2[17:15], tmp2[23:21], tmp2[11:09], tmp2[08:06], tmp2[05:03], tmp2[02:00]} :
                (k3 == 'b100) ? {tmp2[11:09], tmp2[20:18], tmp2[17:15], tmp2[14:12], tmp2[23:21], tmp2[08:06], tmp2[05:03], tmp2[02:00]} :
                (k3 == 'b101) ? {tmp2[08:06], tmp2[20:18], tmp2[17:15], tmp2[14:12], tmp2[11:09], tmp2[23:21], tmp2[05:03], tmp2[02:00]} :
                (k3 == 'b110) ? {tmp2[05:03], tmp2[20:18], tmp2[17:15], tmp2[14:12], tmp2[11:09], tmp2[08:06], tmp2[23:21], tmp2[02:00]} :
                (k3 == 'b111) ? {tmp2[02:00], tmp2[20:18], tmp2[17:15], tmp2[14:12], tmp2[11:09], tmp2[08:06], tmp2[05:03], tmp2[23:21]} :
                                3'bx ;

// number 5
assign k4 = shift_key[11:09];
assign tmp4 =   (k4 == 'b000) ? {tmp3[23:21], tmp3[20:18], tmp3[17:15], tmp3[14:12], tmp3[11:09], tmp3[08:06], tmp3[05:03], tmp3[02:00]} :
                (k4 == 'b001) ? {tmp3[20:18], tmp3[23:21], tmp3[17:15], tmp3[14:12], tmp3[11:09], tmp3[08:06], tmp3[05:03], tmp3[02:00]} :
                (k4 == 'b010) ? {tmp3[17:15], tmp3[20:18], tmp3[23:21], tmp3[14:12], tmp3[11:09], tmp3[08:06], tmp3[05:03], tmp3[02:00]} :
                (k4 == 'b011) ? {tmp3[14:12], tmp3[20:18], tmp3[17:15], tmp3[23:21], tmp3[11:09], tmp3[08:06], tmp3[05:03], tmp3[02:00]} :
                (k4 == 'b100) ? {tmp3[11:09], tmp3[20:18], tmp3[17:15], tmp3[14:12], tmp3[23:21], tmp3[08:06], tmp3[05:03], tmp3[02:00]} :
                (k4 == 'b101) ? {tmp3[08:06], tmp3[20:18], tmp3[17:15], tmp3[14:12], tmp3[11:09], tmp3[23:21], tmp3[05:03], tmp3[02:00]} :
                (k4 == 'b110) ? {tmp3[05:03], tmp3[20:18], tmp3[17:15], tmp3[14:12], tmp3[11:09], tmp3[08:06], tmp3[23:21], tmp3[02:00]} :
                (k4 == 'b111) ? {tmp3[02:00], tmp3[20:18], tmp3[17:15], tmp3[14:12], tmp3[11:09], tmp3[08:06], tmp3[05:03], tmp3[23:21]} :
                                3'bx ;

// number 6
assign k5 = shift_key[08:06];
assign tmp5 =   (k5 == 'b000) ? {tmp4[23:21], tmp4[20:18], tmp4[17:15], tmp4[14:12], tmp4[11:09], tmp4[08:06], tmp4[05:03], tmp4[02:00]} :
                (k5 == 'b001) ? {tmp4[20:18], tmp4[23:21], tmp4[17:15], tmp4[14:12], tmp4[11:09], tmp4[08:06], tmp4[05:03], tmp4[02:00]} :
                (k5 == 'b010) ? {tmp4[17:15], tmp4[20:18], tmp4[23:21], tmp4[14:12], tmp4[11:09], tmp4[08:06], tmp4[05:03], tmp4[02:00]} :
                (k5 == 'b011) ? {tmp4[14:12], tmp4[20:18], tmp4[17:15], tmp4[23:21], tmp4[11:09], tmp4[08:06], tmp4[05:03], tmp4[02:00]} :
                (k5 == 'b100) ? {tmp4[11:09], tmp4[20:18], tmp4[17:15], tmp4[14:12], tmp4[23:21], tmp4[08:06], tmp4[05:03], tmp4[02:00]} :
                (k5 == 'b101) ? {tmp4[08:06], tmp4[20:18], tmp4[17:15], tmp4[14:12], tmp4[11:09], tmp4[23:21], tmp4[05:03], tmp4[02:00]} :
                (k5 == 'b110) ? {tmp4[05:03], tmp4[20:18], tmp4[17:15], tmp4[14:12], tmp4[11:09], tmp4[08:06], tmp4[23:21], tmp4[02:00]} :
                (k5 == 'b111) ? {tmp4[02:00], tmp4[20:18], tmp4[17:15], tmp4[14:12], tmp4[11:09], tmp4[08:06], tmp4[05:03], tmp4[23:21]} :
                                3'bx ;

// number 7
assign k6 = shift_key[05:03];
assign tmp6 =   (k6 == 'b000) ? {tmp5[23:21], tmp5[20:18], tmp5[17:15], tmp5[14:12], tmp5[11:09], tmp5[08:06], tmp5[05:03], tmp5[02:00]} :
                (k6 == 'b001) ? {tmp5[20:18], tmp5[23:21], tmp5[17:15], tmp5[14:12], tmp5[11:09], tmp5[08:06], tmp5[05:03], tmp5[02:00]} :
                (k6 == 'b010) ? {tmp5[17:15], tmp5[20:18], tmp5[23:21], tmp5[14:12], tmp5[11:09], tmp5[08:06], tmp5[05:03], tmp5[02:00]} :
                (k6 == 'b011) ? {tmp5[14:12], tmp5[20:18], tmp5[17:15], tmp5[23:21], tmp5[11:09], tmp5[08:06], tmp5[05:03], tmp5[02:00]} :
                (k6 == 'b100) ? {tmp5[11:09], tmp5[20:18], tmp5[17:15], tmp5[14:12], tmp5[23:21], tmp5[08:06], tmp5[05:03], tmp5[02:00]} :
                (k6 == 'b101) ? {tmp5[08:06], tmp5[20:18], tmp5[17:15], tmp5[14:12], tmp5[11:09], tmp5[23:21], tmp5[05:03], tmp5[02:00]} :
                (k6 == 'b110) ? {tmp5[05:03], tmp5[20:18], tmp5[17:15], tmp5[14:12], tmp5[11:09], tmp5[08:06], tmp5[23:21], tmp5[02:00]} :
                (k6 == 'b111) ? {tmp5[02:00], tmp5[20:18], tmp5[17:15], tmp5[14:12], tmp5[11:09], tmp5[08:06], tmp5[05:03], tmp5[23:21]} :
                                3'bx ;

// number 8
assign k7 = shift_key[02:00];
assign tmp7 =   (k7 == 'b000) ? {tmp6[23:21], tmp6[20:18], tmp6[17:15], tmp6[14:12], tmp6[11:09], tmp6[08:06], tmp6[05:03], tmp6[02:00]} :
                (k7 == 'b001) ? {tmp6[20:18], tmp6[23:21], tmp6[17:15], tmp6[14:12], tmp6[11:09], tmp6[08:06], tmp6[05:03], tmp6[02:00]} :
                (k7 == 'b010) ? {tmp6[17:15], tmp6[20:18], tmp6[23:21], tmp6[14:12], tmp6[11:09], tmp6[08:06], tmp6[05:03], tmp6[02:00]} :
                (k7 == 'b011) ? {tmp6[14:12], tmp6[20:18], tmp6[17:15], tmp6[23:21], tmp6[11:09], tmp6[08:06], tmp6[05:03], tmp6[02:00]} :
                (k7 == 'b100) ? {tmp6[11:09], tmp6[20:18], tmp6[17:15], tmp6[14:12], tmp6[23:21], tmp6[08:06], tmp6[05:03], tmp6[02:00]} :
                (k7 == 'b101) ? {tmp6[08:06], tmp6[20:18], tmp6[17:15], tmp6[14:12], tmp6[11:09], tmp6[23:21], tmp6[05:03], tmp6[02:00]} :
                (k7 == 'b110) ? {tmp6[05:03], tmp6[20:18], tmp6[17:15], tmp6[14:12], tmp6[11:09], tmp6[08:06], tmp6[23:21], tmp6[02:00]} :
                (k7 == 'b111) ? {tmp6[02:00], tmp6[20:18], tmp6[17:15], tmp6[14:12], tmp6[11:09], tmp6[08:06], tmp6[05:03], tmp6[23:21]} :
                                3'bx ;

// final
assign permute_key1 = tmp7;
assign permute_key2 = {
    tmp6[02:00],
    tmp6[05:03],
    tmp6[08:06],
    tmp6[11:09], 
    tmp6[14:12], 
    tmp6[17:15], 
    tmp6[20:18], 
    tmp6[23:21]
    };

endmodule