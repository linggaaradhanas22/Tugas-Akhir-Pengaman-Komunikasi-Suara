library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity lutsin_block is
    Port (
        address      : in  std_logic_vector(9 downto 0);                    -- 640 alamat
        sine_697     : out std_logic_vector(15 downto 0);  
        sine_941     : out std_logic_vector(15 downto 0);  
        sine_1477    : out std_logic_vector(15 downto 0)  
    );
end lutsin_block;

architecture Behavioral of lutsin_block is

    type sample_array is array (0 to 2) of std_logic_vector(15 downto 0);
    type rom_array is array (0 to 639) of sample_array;

    constant rom : rom_array := (
        (x"0000", x"0000", x"0000"), 
        (x"1176", x"1784", x"249A"), 
        (x"2299", x"2E3B", x"4626"), 
        (x"3317", x"435F", x"61D6"), 
        (x"429F", x"5638", x"755A"), 
        (x"50E9", x"6622", x"7F11"), 
        (x"5DB0", x"7292", x"7E2C"), 
        (x"68B5", x"7B1B", x"72BD"), 
        (x"71C6", x"7F73", x"5DB8"), 
        (x"78B6", x"7F75", x"40E0"), 
        (x"7D64", x"7B20", x"1E9D"), 
        (x"7FBA", x"729A", x"F9CB"), 
        (x"7FAC", x"662E", x"D57E"), 
        (x"7D3C", x"5647", x"B4BE"), 
        (x"7873", x"4370", x"9A47"), 
        (x"716A", x"2E4D", x"884F"), 
        (x"6842", x"1797", x"8056"), 
        (x"5D27", x"0013", x"8306"), 
        (x"504E", x"E88F", x"9026"), 
        (x"41F5", x"D1D7", x"A69E"), 
        (x"3260", x"BCB1", x"C48D"), 
        (x"21D9", x"A9D6", x"E773"), 
        (x"10B1", x"99EA", x"0C65"), 
        (x"FF39", x"8D77", x"304F"), 
        (x"EDC4", x"84EA", x"5030"), 
        (x"DCA7", x"808E", x"695F"), 
        (x"CC33", x"8089", x"79C0"), 
        (x"BCB7", x"84DB", x"7FF7"), 
        (x"AE7D", x"8D5D", x"7B7D"), 
        (x"A1C9", x"99C7", x"6CB4"), 
        (x"96D8", x"A9AB", x"54D6"), 
        (x"8DDF", x"BC80", x"35E3"), 
        (x"8708", x"D1A1", x"126F"), 
        (x"8274", x"E856", x"ED71"), 
        (x"803A", x"FFD9", x"CA00"), 
        (x"8063", x"175E", x"AB12"), 
        (x"82EE", x"2E17", x"933B"), 
        (x"87D1", x"433E", x"847A"), 
        (x"8EF3", x"561C", x"800A"), 
        (x"9832", x"660B", x"864A"), 
        (x"A362", x"7280", x"96B4"), 
        (x"B04E", x"7B10", x"AFE9"), 
        (x"BEB7", x"7F70", x"CFCF"), 
        (x"CE58", x"7F79", x"F3BB"), 
        (x"DEE7", x"7B2B", x"18AD"), 
        (x"F015", x"72AB", x"3B90"), 
        (x"018F", x"6645", x"5979"), 
        (x"1301", x"5663", x"6FE9"), 
        (x"2419", x"4390", x"7D01"), 
        (x"3483", x"2E71", x"7FA8"), 
        (x"43F3", x"17BD", x"77A6"), 
        (x"521D", x"003A", x"65A5"), 
        (x"5EBE", x"E8B5", x"4B28"), 
        (x"6999", x"D1FB", x"2A63"), 
        (x"727B", x"BCD2", x"0614"), 
        (x"7938", x"A9F3", x"E144"), 
        (x"7DB2", x"9A01", x"BF04"), 
        (x"7FD2", x"8D88", x"A232"), 
        (x"7F8D", x"84F5", x"8D35"), 
        (x"7CE7", x"8092", x"81CF"), 
        (x"77EA", x"8086", x"80F3"), 
        (x"70AF", x"84D0", x"8AB3"), 
        (x"6759", x"8D4C", x"9E3F"), 
        (x"5C14", x"99B0", x"B9F5"), 
        (x"4F16", x"A98F", x"DB84"), 
        (x"409E", x"BC5F", x"0020"), 
        (x"30F0", x"D17D", x"24B9"), 
        (x"2058", x"E830", x"4641"), 
        (x"0F25", x"FFB3", x"61EB"), 
        (x"FDAA", x"1738", x"7567"), 
        (x"EC3A", x"2DF3", x"7F15"), 
        (x"DB28", x"431E", x"7E26"), 
        (x"CAC7", x"55FF", x"72AE"), 
        (x"BB65", x"65F3", x"5DA2"), 
        (x"AD4B", x"726F", x"40C4"), 
        (x"A0BD", x"7B06", x"1E7E"), 
        (x"95F7", x"7F6C", x"F9AB"), 
        (x"8D2D", x"7F7C", x"D560"), 
        (x"8688", x"7B35", x"B4A4"), 
        (x"8229", x"72BD", x"9A34"), 
        (x"8024", x"665C", x"8843"), 
        (x"8084", x"5680", x"8053"), 
        (x"8346", x"43B1", x"830D"), 
        (x"885C", x"2E95", x"9036"), 
        (x"8FB0", x"17E3", x"A6B5"), 
        (x"991D", x"0061", x"C4A9"), 
        (x"A477", x"E8DB", x"E792"), 
        (x"B187", x"D21F", x"0C85"), 
        (x"C00F", x"BCF3", x"306D"), 
        (x"CFC9", x"AA0F", x"5049"), 
        (x"E069", x"9A18", x"6971"), 
        (x"F1A1", x"8D99", x"79CA"), 
        (x"031E", x"8500", x"7FF8"), 
        (x"148B", x"8096", x"7B75"), 
        (x"2597", x"8082", x"6CA3"), 
        (x"35EE", x"84C6", x"54BE"), 
        (x"4543", x"8D3B", x"35C5"), 
        (x"534D", x"9998", x"124F"), 
        (x"5FC8", x"A972", x"ED51"), 
        (x"6A78", x"BC3E", x"C9E3"), 
        (x"732B", x"D159", x"AAFA"), 
        (x"79B6", x"E80A", x"932A"), 
        (x"7DFB", x"FF8C", x"8472"), 
        (x"7FE4", x"1712", x"800B"), 
        (x"7F6A", x"2DCF", x"8654"), 
        (x"7C8D", x"42FD", x"96C6"), 
        (x"775C", x"55E3", x"B002"), 
        (x"6FF0", x"65DC", x"CFEC"), 
        (x"666C", x"725E", x"F3DB"), 
        (x"5AFD", x"7AFB", x"18CD"), 
        (x"4DDB", x"7F68", x"3BAC"), 
        (x"3F44", x"7F80", x"5990"), 
        (x"2F7E", x"7B40", x"6FF9"), 
        (x"1ED5", x"72CE", x"7D08"), 
        (x"0D99", x"6673", x"7FA6"), 
        (x"FC1B", x"569C", x"779A"), 
        (x"EAB0", x"43D2", x"6592"), 
        (x"D9AB", x"2EB9", x"4B0E"), 
        (x"C95D", x"1809", x"2A45"), 
        (x"BA15", x"0087", x"05F4"), 
        (x"AC1C", x"E901", x"E124"), 
        (x"9FB4", x"D243", x"BEE8"), 
        (x"9519", x"BD14", x"A21C"), 
        (x"8C7F", x"AA2C", x"8D27"), 
        (x"860D", x"9A30", x"81C9"), 
        (x"81E2", x"8DAB", x"80F6"), 
        (x"8014", x"850A", x"8AC0"), 
        (x"80AA", x"8099", x"9E53"), 
        (x"83A2", x"807F", x"BA10"), 
        (x"88ED", x"84BB", x"DBA3"), 
        (x"9072", x"8D2A", x"0040"), 
        (x"9A0D", x"9981", x"24D8"), 
        (x"A590", x"A956", x"465C"), 
        (x"B2C4", x"BC1E", x"61FF"), 
        (x"C16A", x"D135", x"7574"), 
        (x"D13B", x"E7E4", x"7F19"), 
        (x"E1EC", x"FF66", x"7E21"), 
        (x"F32E", x"16EC", x"72A0"), 
        (x"04AC", x"2DAB", x"5D8C"), 
        (x"1615", x"42DC", x"40A9"), 
        (x"2713", x"55C6", x"1E5F"), 
        (x"3757", x"65C5", x"F98B"), 
        (x"4692", x"724C", x"D542"), 
        (x"547A", x"7AF0", x"B48A"), 
        (x"60CF", x"7F65", x"9A20"), 
        (x"6B54", x"7F83", x"8838"), 
        (x"73D7", x"7B4A", x"8051"), 
        (x"7A2F", x"72DF", x"8314"), 
        (x"7E3F", x"668A", x"9045"), 
        (x"7FF2", x"56B8", x"A6CC"), 
        (x"7F41", x"43F3", x"C4C6"), 
        (x"7C2F", x"2EDD", x"E7B2"), 
        (x"76CA", x"182F", x"0CA5"), 
        (x"6F2C", x"00AE", x"308B"), 
        (x"657A", x"E927", x"5062"), 
        (x"59E3", x"D267", x"6983"), 
        (x"4C9D", x"BD35", x"79D4"), 
        (x"3DE8", x"AA48", x"7FF8"), 
        (x"2E0B", x"9A47", x"7B6C"), 
        (x"1D52", x"8DBC", x"6C92"), 
        (x"0C0C", x"8515", x"54A6"), 
        (x"FA8C", x"809D", x"35A8"), 
        (x"E927", x"807B", x"122F"), 
        (x"D82F", x"84B1", x"ED32"), 
        (x"C7F5", x"8D19", x"C9C6"), 
        (x"B8C8", x"996A", x"AAE2"), 
        (x"AAF0", x"A939", x"9319"), 
        (x"9EAF", x"BBFD", x"8469"), 
        (x"9440", x"D111", x"800C"), 
        (x"8BD5", x"E7BE", x"865E"), 
        (x"8596", x"FF3F", x"96D8"), 
        (x"81A1", x"16C6", x"B01B"), 
        (x"8008", x"2D87", x"D00A"), 
        (x"80D5", x"42BB", x"F3FB"), 
        (x"8402", x"55A9", x"18EC"), 
        (x"8981", x"65AD", x"3BC9"), 
        (x"9137", x"723B", x"59A7"), 
        (x"9B00", x"7AE6", x"7009"), 
        (x"A6AC", x"7F61", x"7D0F"), 
        (x"B403", x"7F86", x"7FA3"), 
        (x"C2C7", x"7B54", x"778F"), 
        (x"D2AF", x"72F0", x"657E"), 
        (x"E371", x"66A1", x"4AF4"), 
        (x"F4BB", x"56D5", x"2A26"), 
        (x"063B", x"4413", x"05D4"), 
        (x"179D", x"2F01", x"E105"), 
        (x"288F", x"1855", x"BECD"), 
        (x"38BE", x"00D4", x"A206"), 
        (x"47DD", x"E94D", x"8D19"), 
        (x"55A4", x"D28B", x"81C4"), 
        (x"61D2", x"BD56", x"80FA"), 
        (x"6C2B", x"AA65", x"8ACC"), 
        (x"747E", x"9A5F", x"9E68"), 
        (x"7AA4", x"8DCE", x"BA2B"), 
        (x"7E7E", x"8520", x"DBC2"), 
        (x"7FFB", x"80A1", x"0061"), 
        (x"7F14", x"8078", x"24F7"), 
        (x"7BCC", x"84A6", x"4677"), 
        (x"7633", x"8D08", x"6214"), 
        (x"6E64", x"9953", x"7581"), 
        (x"6485", x"A91D", x"7F1D"), 
        (x"58C5", x"BBDC", x"7E1B"), 
        (x"4B5C", x"D0ED", x"7292"), 
        (x"3C8A", x"E798", x"5D76"), 
        (x"2C96", x"FF18", x"408D"), 
        (x"1BCD", x"16A0", x"1E3F"), 
        (x"0A7E", x"2D63", x"F96B"), 
        (x"F8FE", x"429A", x"D523"), 
        (x"E79F", x"558D", x"B470"), 
        (x"D6B4", x"6596", x"9A0D"), 
        (x"C690", x"722A", x"882D"), 
        (x"B77E", x"7ADB", x"804F"), 
        (x"A9C8", x"7F5D", x"831B"), 
        (x"9DAE", x"7F8A", x"9055"), 
        (x"936B", x"7B5F", x"A6E3"), 
        (x"8B30", x"7301", x"C4E2"), 
        (x"8523", x"66B8", x"E7D1"), 
        (x"8164", x"56F1", x"0CC5"), 
        (x"8002", x"4434", x"30A9"), 
        (x"8105", x"2F25", x"507B"), 
        (x"8468", x"187A", x"6995"), 
        (x"8A1A", x"00FB", x"79DE"), 
        (x"9201", x"E973", x"7FF9"), 
        (x"9BF7", x"D2AF", x"7B64"), 
        (x"A7CB", x"BD77", x"6C81"), 
        (x"B546", x"AA82", x"548E"), 
        (x"C426", x"9A76", x"358B"), 
        (x"D425", x"8DDF", x"120F"), 
        (x"E4F6", x"852B", x"ED12"), 
        (x"F648", x"80A5", x"C9A9"), 
        (x"07C9", x"8075", x"AACA"), 
        (x"1925", x"849C", x"9308"), 
        (x"2A08", x"8CF7", x"8461"), 
        (x"3A22", x"993C", x"800D"), 
        (x"4926", x"A901", x"8668"), 
        (x"56CB", x"BBBC", x"96EB"), 
        (x"62D1", x"D0C9", x"B034"), 
        (x"6CFE", x"E773", x"D028"), 
        (x"7521", x"FEF2", x"F41B"), 
        (x"7B14", x"167A", x"190C"), 
        (x"7EB9", x"2D3F", x"3BE5"), 
        (x"7FFF", x"4279", x"59BE"), 
        (x"7EE1", x"5570", x"7018"), 
        (x"7B64", x"657E", x"7D16"), 
        (x"7598", x"7218", x"7FA1"), 
        (x"6D98", x"7AD0", x"7783"), 
        (x"638C", x"7F59", x"656B"), 
        (x"57A4", x"7F8D", x"4ADA"), 
        (x"4A18", x"7B69", x"2A08"), 
        (x"3B29", x"7312", x"05B4"), 
        (x"2B1F", x"66D0", x"E0E6"), 
        (x"1A47", x"570D", x"BEB1"), 
        (x"08F1", x"4455", x"A1F0"), 
        (x"F770", x"2F49", x"8D0B"), 
        (x"E618", x"18A0", x"81BF"), 
        (x"D53C", x"0122", x"80FE"), 
        (x"C52C", x"E999", x"8AD9"), 
        (x"B637", x"D2D3", x"9E7D"), 
        (x"A8A3", x"BD98", x"BA46"), 
        (x"9CB0", x"AA9F", x"DBE1"), 
        (x"929A", x"9A8E", x"0081"), 
        (x"8A8F", x"8DF1", x"2516"), 
        (x"84B6", x"8536", x"4692"), 
        (x"812B", x"80A9", x"6229"), 
        (x"8000", x"8071", x"758D"), 
        (x"8139", x"8492", x"7F21"), 
        (x"84D2", x"8CE6", x"7E16"), 
        (x"8AB8", x"9925", x"7283"), 
        (x"92CF", x"A8E4", x"5D60"), 
        (x"9CF1", x"BB9B", x"4071"), 
        (x"A8EE", x"D0A5", x"1E20"), 
        (x"B68B", x"E74D", x"F94B"), 
        (x"C588", x"FECB", x"D505"), 
        (x"D59D", x"1654", x"B456"), 
        (x"E67D", x"2D1B", x"99F9"), 
        (x"F7D6", x"4258", x"8821"), 
        (x"0957", x"5553", x"804C"), 
        (x"1AAC", x"6567", x"8322"), 
        (x"2B80", x"7207", x"9065"), 
        (x"3B84", x"7AC5", x"A6FA"), 
        (x"4A6C", x"7F55", x"C4FF"), 
        (x"57EF", x"7F90", x"E7F1"), 
        (x"63CD", x"7B73", x"0CE5"), 
        (x"6DCD", x"7323", x"30C6"), 
        (x"75C0", x"66E6", x"5094"), 
        (x"7B7F", x"572A", x"69A7"), 
        (x"7EEF", x"4475", x"79E8"), 
        (x"7FFF", x"2F6C", x"7FFA"), 
        (x"7EAA", x"18C6", x"7B5B"), 
        (x"7AF7", x"0148", x"6C70"), 
        (x"74F8", x"E9BF", x"5476"), 
        (x"6CC8", x"D2F8", x"356E"), 
        (x"6290", x"BDB9", x"11F0"), 
        (x"5680", x"AABB", x"ECF2"), 
        (x"48D1", x"9AA5", x"C98C"), 
        (x"39C6", x"8E02", x"AAB2"), 
        (x"29A7", x"8541", x"92F8"), 
        (x"18C0", x"80AD", x"8459"), 
        (x"0763", x"806E", x"800D"), 
        (x"F5E2", x"8488", x"8672"), 
        (x"E492", x"8CD5", x"96FD"), 
        (x"D3C5", x"990E", x"B04E"), 
        (x"C3CB", x"A8C8", x"D046"), 
        (x"B4F2", x"BB7A", x"F43B"), 
        (x"A781", x"D082", x"192B"), 
        (x"9BB7", x"E727", x"3C02"), 
        (x"91CD", x"FEA5", x"59D5"), 
        (x"89F2", x"162E", x"7028"), 
        (x"844D", x"2CF6", x"7D1D"), 
        (x"80F8", x"4237", x"7F9E"), 
        (x"8003", x"5536", x"7778"), 
        (x"8173", x"654F", x"6557"), 
        (x"8541", x"71F5", x"4ABF"), 
        (x"8B5A", x"7ABA", x"29EA"), 
        (x"93A1", x"7F51", x"0594"), 
        (x"9DF0", x"7F93", x"E0C7"), 
        (x"AA14", x"7B7D", x"BE95"), 
        (x"B7D3", x"7333", x"A1DA"), 
        (x"C6EC", x"66FD", x"8CFC"), 
        (x"D716", x"5746", x"81BA"), 
        (x"E804", x"4496", x"8102"), 
        (x"F965", x"2F90", x"8AE6"), 
        (x"0AE5", x"18EC", x"9E92"), 
        (x"1C31", x"016F", x"BA61"), 
        (x"2CF6", x"E9E5", x"DC00"), 
        (x"3CE4", x"D31C", x"00A1"), 
        (x"4BAF", x"BDDA", x"2534"), 
        (x"590F", x"AAD8", x"46AC"), 
        (x"64C5", x"9ABD", x"623D"), 
        (x"6E98", x"8E14", x"759A"), 
        (x"765A", x"854B", x"7F24"), 
        (x"7BE6", x"80B1", x"7E10"), 
        (x"7F20", x"806B", x"7275"), 
        (x"7FFA", x"847E", x"5D4A"), 
        (x"7E6F", x"8CC4", x"4055"), 
        (x"7A86", x"98F7", x"1E01"), 
        (x"7454", x"A8AC", x"F92B"), 
        (x"6BF4", x"BB5A", x"D4E7"), 
        (x"618F", x"D05E", x"B43C"), 
        (x"5558", x"E701", x"99E6"), 
        (x"4788", x"FE7E", x"8816"), 
        (x"3861", x"1608", x"804A"), 
        (x"282D", x"2CD2", x"8329"), 
        (x"1738", x"4216", x"9075"), 
        (x"05D4", x"5519", x"A711"), 
        (x"F454", x"6538", x"C51B"), 
        (x"E30C", x"71E3", x"E811"), 
        (x"D24F", x"7AAF", x"0D05"), 
        (x"C26C", x"7F4D", x"30E4"), 
        (x"B3B1", x"7F96", x"50AD"), 
        (x"A662", x"7B88", x"69BA"), 
        (x"9AC1", x"7344", x"79F1"), 
        (x"9104", x"6714", x"7FFA"), 
        (x"895A", x"5762", x"7B53"), 
        (x"83E9", x"44B7", x"6C5F"), 
        (x"80C9", x"2FB4", x"545D"), 
        (x"800B", x"1912", x"3550"), 
        (x"81B1", x"0195", x"11D0"), 
        (x"85B4", x"EA0B", x"ECD2"), 
        (x"8C00", x"D340", x"C96F"), 
        (x"9478", x"BDFB", x"AA9A"), 
        (x"9EF2", x"AAF5", x"92E7"), 
        (x"AB3D", x"9AD4", x"8450"), 
        (x"B91E", x"8E25", x"800E"), 
        (x"C852", x"8557", x"867C"), 
        (x"D891", x"80B5", x"970F"), 
        (x"E98C", x"8068", x"B067"), 
        (x"FAF3", x"8473", x"D064"), 
        (x"0C72", x"8CB3", x"F45B"), 
        (x"1DB6", x"98E0", x"194B"), 
        (x"2E6B", x"A890", x"3C1E"), 
        (x"3E42", x"BB39", x"59EC"), 
        (x"4CEF", x"D03A", x"7037"), 
        (x"5A2C", x"E6DB", x"7D23"), 
        (x"65B9", x"FE57", x"7F9C"), 
        (x"6F5F", x"15E2", x"776C"), 
        (x"76F0", x"2CAE", x"6543"), 
        (x"7C47", x"41F5", x"4AA5"), 
        (x"7F4C", x"54FD", x"29CB"), 
        (x"7FEF", x"6520", x"0574"), 
        (x"7E2E", x"71D2", x"E0A8"), 
        (x"7A11", x"7AA4", x"BE7A"), 
        (x"73AB", x"7F49", x"A1C5"), 
        (x"6B1B", x"7F99", x"8CEE"), 
        (x"608B", x"7B92", x"81B4"), 
        (x"542D", x"7355", x"8106"), 
        (x"463C", x"672B", x"8AF3"), 
        (x"36FA", x"577E", x"9EA7"), 
        (x"26B1", x"44D7", x"BA7C"), 
        (x"15AF", x"2FD8", x"DC1F"), 
        (x"0446", x"1938", x"00C1"), 
        (x"F2C7", x"01BC", x"2553"), 
        (x"E188", x"EA31", x"46C7"), 
        (x"D0DB", x"D364", x"6252"), 
        (x"C110", x"BE1C", x"75A7"), 
        (x"B272", x"AB12", x"7F28"), 
        (x"A547", x"9AEC", x"7E0B"), 
        (x"99CE", x"8E37", x"7267"), 
        (x"903F", x"8562", x"5D34"), 
        (x"88C7", x"80B9", x"403A"), 
        (x"8389", x"8065", x"1DE2"), 
        (x"80A0", x"8469", x"F90B"), 
        (x"8018", x"8CA3", x"D4C9"), 
        (x"81F4", x"98C9", x"B422"), 
        (x"862C", x"A874", x"99D2"), 
        (x"8CAB", x"BB19", x"880B"), 
        (x"9552", x"D016", x"8048"), 
        (x"9FF8", x"E6B5", x"8330"), 
        (x"AC6A", x"FE31", x"9084"), 
        (x"BA6B", x"15BC", x"A728"), 
        (x"C9BA", x"2C8A", x"C538"), 
        (x"DA0D", x"41D4", x"E830"), 
        (x"EB15", x"54E0", x"0D25"), 
        (x"FC82", x"6508", x"3102"), 
        (x"0DFF", x"71C0", x"50C6"), 
        (x"1F39", x"7A99", x"69CC"), 
        (x"2FDE", x"7F45", x"79FB"), 
        (x"3F9D", x"7F9C", x"7FFB"), 
        (x"4E2C", x"7B9C", x"7B4A"), 
        (x"5B45", x"7366", x"6C4D"), 
        (x"66A9", x"6742", x"5445"), 
        (x"7022", x"579B", x"3533"), 
        (x"7781", x"44F8", x"11B0"), 
        (x"7CA5", x"2FFC", x"ECB2"), 
        (x"7F73", x"195E", x"C952"), 
        (x"7FE0", x"01E3", x"AA82"), 
        (x"7DE9", x"EA57", x"92D6"), 
        (x"7996", x"D388", x"8448"), 
        (x"72FE", x"BE3D", x"800F"), 
        (x"6A3F", x"AB2F", x"8686"), 
        (x"5F84", x"9B04", x"9722"), 
        (x"52FF", x"8E49", x"B080"), 
        (x"44ED", x"856D", x"D082"), 
        (x"3591", x"80BD", x"F47B"), 
        (x"2534", x"8062", x"196A"), 
        (x"1426", x"845F", x"3C3A"), 
        (x"02B7", x"8C92", x"5A03"), 
        (x"F13B", x"98B3", x"7047"), 
        (x"E006", x"A857", x"7D2A"), 
        (x"CF69", x"BAF8", x"7F99"), 
        (x"BFB6", x"CFF2", x"7761"), 
        (x"B136", x"E68F", x"6530"), 
        (x"A42F", x"FE0A", x"4A8B"), 
        (x"98E0", x"1596", x"29AD"), 
        (x"8F7F", x"2C66", x"0554"), 
        (x"8838", x"41B3", x"E088"), 
        (x"832F", x"54C3", x"BE5E"), 
        (x"807B", x"64F0", x"A1AF"), 
        (x"8029", x"71AE", x"8CE0"), 
        (x"823C", x"7A8E", x"81AF"), 
        (x"86A9", x"7F41", x"810B"), 
        (x"8D5A", x"7F9F", x"8B00"), 
        (x"9631", x"7BA6", x"9EBC"), 
        (x"A102", x"7376", x"BA97"), 
        (x"AD99", x"6759", x"DC3E"), 
        (x"BBBC", x"57B7", x"00E1"), 
        (x"CB25", x"4518", x"2572"), 
        (x"DB8B", x"3020", x"46E2"), 
        (x"EC9F", x"1983", x"6267"), 
        (x"FE11", x"0209", x"75B3"), 
        (x"0F8B", x"EA7D", x"7F2C"), 
        (x"20BB", x"D3AC", x"7E05"), 
        (x"314F", x"BE5E", x"7258"), 
        (x"40F6", x"AB4C", x"5D1E"), 
        (x"4F67", x"9B1B", x"401E"), 
        (x"5C5B", x"8E5A", x"1DC2"), 
        (x"6795", x"8578", x"F8EB"), 
        (x"70E0", x"80C1", x"D4AA"), 
        (x"780E", x"805F", x"B409"), 
        (x"7CFD", x"8455", x"99BF"), 
        (x"7F96", x"8C81", x"8800"), 
        (x"7FCC", x"989C", x"8046"), 
        (x"7D9E", x"A83B", x"8337"), 
        (x"7917", x"BAD8", x"9094"), 
        (x"724C", x"CFCF", x"A740"), 
        (x"695F", x"E66A", x"C555"), 
        (x"5E78", x"FDE4", x"E850"), 
        (x"51CE", x"1570", x"0D45"), 
        (x"439B", x"2C41", x"311F"), 
        (x"3425", x"4191", x"50DF"), 
        (x"23B6", x"54A6", x"69DE"), 
        (x"129C", x"64D9", x"7A05"), 
        (x"0128", x"719D", x"7FFB"), 
        (x"EFAF", x"7A83", x"7B41"), 
        (x"DE84", x"7F3D", x"6C3C"), 
        (x"CDF9", x"7FA2", x"542D"), 
        (x"BE5E", x"7BB0", x"3516"), 
        (x"AFFD", x"7387", x"1190"), 
        (x"A31B", x"6770", x"EC93"), 
        (x"97F6", x"57D3", x"C934"), 
        (x"8EC3", x"4539", x"AA6A"), 
        (x"87AE", x"3043", x"92C5"), 
        (x"82D9", x"19A9", x"8440"), 
        (x"805B", x"0230", x"8010"), 
        (x"8040", x"EAA3", x"8690"), 
        (x"8289", x"D3D1", x"9734"), 
        (x"872A", x"BE7F", x"B099"), 
        (x"8E0E", x"AB69", x"D0A0"), 
        (x"9713", x"9B33", x"F49B"), 
        (x"A20F", x"8E6C", x"198A"), 
        (x"AECC", x"8583", x"3C57"), 
        (x"BD0E", x"80C5", x"5A1A"), 
        (x"CC91", x"805C", x"7056"), 
        (x"DD0A", x"844B", x"7D31"), 
        (x"EE2A", x"8C71", x"7F97"), 
        (x"FF9F", x"9885", x"7755"), 
        (x"1117", x"A81F", x"651C"), 
        (x"223C", x"BAB7", x"4A71"), 
        (x"32BE", x"CFAB", x"298E"), 
        (x"424D", x"E644", x"0533"), 
        (x"509E", x"FDBD", x"E069"), 
        (x"5D6E", x"154A", x"BE42"), 
        (x"687E", x"2C1D", x"A199"), 
        (x"719A", x"4170", x"8CD2"), 
        (x"7896", x"5489", x"81AA"), 
        (x"7D51", x"64C1", x"810F"), 
        (x"7FB4", x"718B", x"8B0D"), 
        (x"7FB3", x"7A77", x"9ED1"), 
        (x"7D4F", x"7F39", x"BAB2"), 
        (x"7894", x"7FA5", x"DC5D"), 
        (x"7197", x"7BBA", x"0101"), 
        (x"687A", x"7398", x"2591"), 
        (x"5D69", x"6786", x"46FD"), 
        (x"5099", x"57EF", x"627B"), 
        (x"4247", x"4559", x"75C0"), 
        (x"32B8", x"3067", x"7F2F"), 
        (x"2236", x"19CF", x"7DFF"), 
        (x"1110", x"0256", x"724A"), 
        (x"FF99", x"EAC9", x"5D08"), 
        (x"EE24", x"D3F5", x"4002"), 
        (x"DD04", x"BEA0", x"1DA3"), 
        (x"CC8B", x"AB86", x"F8CA"), 
        (x"BD09", x"9B4B", x"D48C"), 
        (x"AEC7", x"8E7E", x"B3EF"), 
        (x"A20A", x"858E", x"99AC"), 
        (x"970F", x"80C9", x"87F4"), 
        (x"8E0B", x"8059", x"8044"), 
        (x"8728", x"8442", x"833E"), 
        (x"8287", x"8C60", x"90A4"), 
        (x"803F", x"986E", x"A757"), 
        (x"805B", x"A803", x"C571"), 
        (x"82DA", x"BA97", x"E86F"), 
        (x"87B0", x"CF87", x"0D65"), 
        (x"8EC6", x"E61E", x"313D"), 
        (x"97FA", x"FD96", x"50F8"), 
        (x"A320", x"1524", x"69F0"), 
        (x"B002", x"2BF9", x"7A0F"), 
        (x"BE64", x"414F", x"7FFC"), 
        (x"CDFF", x"546C", x"7B39"), 
        (x"DE8A", x"64A9", x"6C2B"), 
        (x"EFB5", x"7179", x"5415"), 
        (x"012E", x"7A6C", x"34F9"), 
        (x"12A2", x"7F34", x"1170"), 
        (x"23BC", x"7FA8", x"EC73"), 
        (x"342B", x"7BC3", x"C917"), 
        (x"43A1", x"73A8", x"AA52"), 
        (x"51D3", x"679D", x"92B4"), 
        (x"5E7D", x"580B", x"8438"), 
        (x"6962", x"457A", x"8011"), 
        (x"724F", x"308B", x"869A"), 
        (x"7919", x"19F5", x"9747"), 
        (x"7DA0", x"027D", x"B0B2"), 
        (x"7FCC", x"EAEF", x"D0BD"), 
        (x"7F95", x"D419", x"F4BB"), 
        (x"7CFC", x"BEC2", x"19A9"), 
        (x"780C", x"ABA3", x"3C73"), 
        (x"70DD", x"9B63", x"5A30"), 
        (x"6792", x"8E90", x"7066"), 
        (x"5C57", x"8599", x"7D38"), 
        (x"4F62", x"80CE", x"7F94"), 
        (x"40F1", x"8056", x"7749"), 
        (x"3149", x"8438", x"6508"), 
        (x"20B5", x"8C50", x"4A57"), 
        (x"0F85", x"9858", x"2970"), 
        (x"FE0A", x"A7E7", x"0513"), 
        (x"EC99", x"BA76", x"E04A"), 
        (x"DB84", x"CF63", x"BE27"), 
        (x"CB1F", x"E5F8", x"A183"), 
        (x"BBB6", x"FD70", x"8CC4"), 
        (x"AD94", x"14FE", x"81A5"), 
        (x"A0FD", x"2BD5", x"8113"), 
        (x"962D", x"412E", x"8B1B"), 
        (x"8D57", x"544F", x"9EE6"), 
        (x"86A7", x"6491", x"BACD"), 
        (x"823B", x"7167", x"DC7B"), 
        (x"8029", x"7A61", x"0122"), 
        (x"807B", x"7F30", x"25AF"), 
        (x"8330", x"7FAB", x"4718"), 
        (x"883A", x"7BCD", x"6290"), 
        (x"8F82", x"73B9", x"75CD"), 
        (x"98E4", x"67B4", x"7F33"), 
        (x"A434", x"5827", x"7DFA"), 
        (x"B13B", x"459A", x"723B"), 
        (x"BFBB", x"30AE", x"5CF2"), 
        (x"CF6F", x"1A1B", x"3FE6"), 
        (x"E00C", x"02A4", x"1D84"), 
        (x"F141", x"EB15", x"F8AA"), 
        (x"02BD", x"D43D", x"D46E"), 
        (x"142C", x"BEE3", x"B3D5"), 
        (x"253B", x"ABC0", x"9998"), 
        (x"3597", x"9B7B", x"87E9"), 
        (x"44F2", x"8EA2", x"8042"), 
        (x"5304", x"85A5", x"8346"), 
        (x"5F88", x"80D2", x"90B4"), 
        (x"6A43", x"8054", x"A76E"), 
        (x"7301", x"842E", x"C58E"), 
        (x"7998", x"8C3F", x"E88F"), 
        (x"7DEA", x"9841", x"0D85"), 
        (x"7FE0", x"A7CB", x"315B"), 
        (x"7F73", x"BA56", x"5111"), 
        (x"7CA3", x"CF40", x"6A02"), 
        (x"777F", x"E5D2", x"7A18"), 
        (x"701E", x"FD49", x"7FFC"), 
        (x"66A5", x"14D8", x"7B30"), 
        (x"5B41", x"2BB0", x"6C1A"), 
        (x"4E27", x"410D", x"53FC"), 
        (x"3F98", x"5432", x"34DB"), 
        (x"2FD8", x"6479", x"1150"), 
        (x"1F33", x"7155", x"EC53"), 
        (x"0DF9", x"7A56", x"C8FA"), 
        (x"FC7B", x"7F2C", x"AA3A"), 
        (x"EB0F", x"7FAE", x"92A4"), 
        (x"DA07", x"7BD7", x"842F"), 
        (x"C9B4", x"73C9", x"8012"), 
        (x"BA66", x"67CA", x"86A5"), 
        (x"AC65", x"5843", x"9759"), 
        (x"9FF4", x"45BA", x"B0CC"), 
        (x"954F", x"30D2", x"D0DB"), 
        (x"8CA8", x"1A41", x"F4DB"), 
        (x"862A", x"02CA", x"19C9"), 
        (x"81F3", x"EB3B", x"3C8F"), 
        (x"8018", x"D462", x"5A47"), 
        (x"80A0", x"BF04", x"7075"), 
        (x"838B", x"ABDD", x"7D3E"), 
        (x"88C9", x"9B93", x"7F92"), 
        (x"9042", x"8EB4", x"773E"), 
        (x"99D2", x"85B0", x"64F4"), 
        (x"A54C", x"80D6", x"4A3D"), 
        (x"B277", x"8051", x"2952"), 
        (x"C116", x"8424", x"04F3")
    );

begin
    sine_697   <= rom(to_integer(unsigned(address)))(0);
    sine_941   <= rom(to_integer(unsigned(address)))(1);
    sine_1477  <= rom(to_integer(unsigned(address)))(2);
end Behavioral;
