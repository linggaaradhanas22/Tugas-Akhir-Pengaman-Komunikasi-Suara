
// module for complex multiplication
// for WIDTH = 16, works with frac=15 

module Multiply #(
    parameter   WIDTH = 16
)(
    input   signed  [WIDTH-1:0] a_re,
    input   signed  [WIDTH-1:0] a_im,
    input   signed  [WIDTH-1:0] b_re,
    input   signed  [WIDTH-1:0] b_im,

    output  signed  [WIDTH-1:0] m_re,
    output  signed  [WIDTH-1:0] m_im
);

wire signed [WIDTH*2-1:0]   arbr, arbi, aibr, aibi;
wire signed [WIDTH-1:0]     sc_arbr, sc_arbi, sc_aibr, sc_aibi;

//  signed multiplication
assign  arbr = a_re * b_re;
assign  arbi = a_re * b_im;
assign  aibr = a_im * b_re;
assign  aibi = a_im * b_im;

//  scaling
assign  sc_arbr = arbr >>> (WIDTH - 1);
assign  sc_arbi = arbi >>> (WIDTH - 1);
assign  sc_aibr = aibr >>> (WIDTH - 1);
assign  sc_aibi = aibi >>> (WIDTH - 1);

//  sub/add
//  sub/add may overflow if unnormalized data is input
assign  m_re = sc_arbr - sc_aibi;
assign  m_im = sc_arbi + sc_aibr;

endmodule